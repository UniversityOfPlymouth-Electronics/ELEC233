library verilog;
use verilog.vl_types.all;
entity behavioural_vlg_check_tst is
    port(
        Y_behave        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end behavioural_vlg_check_tst;
