library verilog;
use verilog.vl_types.all;
entity behavioural_vlg_vec_tst is
end behavioural_vlg_vec_tst;
